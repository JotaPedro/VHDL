----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    20:02:08 04/16/2016 
-- Design Name: 
-- Module Name:    FullSub - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity FullSub is
    Port ( Ax : in  STD_LOGIC;
           Bx : in  STD_LOGIC;
           Bw_in : in  STD_LOGIC;
           Result : out  STD_LOGIC;
           Bw_out : out  STD_LOGIC);
end FullSub;

architecture Behavioral of FullSub is

begin


end Behavioral;

